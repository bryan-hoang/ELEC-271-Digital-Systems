library ieee;
use ieee.std_logic_1164.all;

package my_components is -- Declares custom components found in other files

component lab5
  port (
        -- Fill in the port definitions
        -- as in the entity VHDL file
       );
end component;

component fsm
  port (
        -- Fill in the port definitions
        -- as in the entity VHDL file
       );
end component;

end package;
